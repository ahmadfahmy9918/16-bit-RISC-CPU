LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RED IS
PORT(
	RED_in : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	RED_out: OUT UNSIGNED(7 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE Behavior OF RED IS 
BEGIN
	RED_out <= UNSIGNED(RED_IN(7 DOWNTO 0));
END Behavior;